library verilog;
use verilog.vl_types.all;
entity ej1labfpga_vlg_vec_tst is
end ej1labfpga_vlg_vec_tst;
