library verilog;
use verilog.vl_types.all;
entity Estados_vlg_vec_tst is
end Estados_vlg_vec_tst;
