library verilog;
use verilog.vl_types.all;
entity esquematicoC_vlg_check_tst is
    port(
        borrout         : in     vl_logic;
        r1              : in     vl_logic;
        r2              : in     vl_logic;
        r3              : in     vl_logic;
        r4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end esquematicoC_vlg_check_tst;
