library verilog;
use verilog.vl_types.all;
entity esclavo_vlg_vec_tst is
end esclavo_vlg_vec_tst;
