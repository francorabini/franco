library verilog;
use verilog.vl_types.all;
entity restador_vlg_vec_tst is
end restador_vlg_vec_tst;
