library verilog;
use verilog.vl_types.all;
entity esquematicoC_vlg_vec_tst is
end esquematicoC_vlg_vec_tst;
