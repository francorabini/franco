library IEEE;
use IEEE.STD_LOGIC_1164.ALL 
entity ej1labfpga is 
port ( SW1 : in STD_LOGIC;
SW2 : in STD_LOGIC;
SW3 : in STD_lOGIC;
LED : out STD_LOGIC);
end ej1labfpga;

